`timescale 1ns / 1ps

module Temporizer(
    input clk,
    input upBottom,
    input downButton,
    input LeftButton,
    input RightButton,
    input actionButton,
    output _time,
    output state
    );







endmodule
