`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:28:42 09/01/2016 
// Design Name: 
// Module Name:    VideoMemorie 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module VideoMemorie(
    input [11:0] Bitscolores,
    input Cordanadas,
    input Pxcount,
    output Vr,
    output Vb,
    output Vg
    );


endmodule
